** sch_path: /home/ilker/Projects/OpenICEDA/Project/xschem/amplifier.sch
**.subckt amplifier Vin Vin out
*.ipin Vin
*.ipin Vin
*.opin out
Vin Vin GND pulse(0 0.1 1ns 1ns 1n 4ns 10ns)
V1 VDD GND 1.8
XM1 out Vin net1 VDD sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
R1 VDD Vin 1k m=1
R2 Vin GND 1k m=1
R3 VDD out 1k m=1
R4 net1 GND 200 m=1
**** begin user architecture code

** opencircuitdesign pdks install
.lib /home/ilker/Projects/OpenICEDA/src/open_pdks/sky130/sky130A/libs.tech/ngspice/sky130.lib.spice tt



.tran 0.01n 1u
.save all


**** end user architecture code
**.ends
.GLOBAL VDD
.GLOBAL GND
.end
