** sch_path: /home/ilker/Projects/OpenICEDA/Project/xschem/untitled-1.sch
**.subckt untitled-1 Vin Vin out
*.ipin Vin
*.ipin Vin
*.opin out
XM2 out Vin GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=5 m=5
Vin Vin GND SIN(-200m 200m 2000000 0 0)
vcc VDD GND 1.8
R1 VDD out 200k m=1
Vin3 __UNCONNECTED_PIN__0 __UNCONNECTED_PIN__1 pulse(-200m 200m 1ns 1ns 1ns 50ns 100ns)
**** begin user architecture code

* this option enables mos model bin
* selection based on W/NF instead of W
.option wnflag=1
*.option savecurrents
.control
tran 0.01n 1us
plot v(vg) vs v(vd)
plot v(vg) vs v(vvs)
plot v(vvs) vs v(vd)
plot v(out) v(vg)
plot v(Vin) vs v(out)
plot all.vcc#branch vs v(Vin)
plot all.vcc#branch vs v(out)
op
.endc



** opencircuitdesign pdks install
.lib /home/ilker/Projects/OpenICEDA/src/open_pdks/sky130/sky130A/libs.tech/ngspice/sky130.lib.spice tt


**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.end
