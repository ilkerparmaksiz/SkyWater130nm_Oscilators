** sch_path: /home/ilker/Projects/OpenICEDA/Project/xschem/untitled-2.sch
**.subckt untitled-2 vdd vdd vdd in in out
*.ipin vdd
*.ipin vdd
*.ipin vdd
*.ipin in
*.ipin in
*.opin out
XQ1 net2 net1 net3 sky130_fd_pr__pnp_05v5_W3p40L3p40
R1 net1 vdd 22k m=1
R2 GND net2 5.1k m=1
R3 GND net1 90k m=1
R4 net3 vdd 1.2k m=1
C1 in net1 10u m=1
V1 vdd GND 15
C2 net2 out 100u m=1
V2 in GND SIN(0 100m 10000 0 0)
R5 GND out 1k m=1
**** begin user architecture code

** opencircuitdesign pdks install
.lib /home/ilker/Projects/OpenICEDA/src/open_pdks/sky130/sky130A/libs.tech/ngspice/sky130.lib.spice tt



* this option enables mos model bin
* selection based on W/NF instead of W
.option wnflag=1
*.option savecurrents
.control
tran 1us 1m
plot v(in) v(out)
op
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
