** sch_path: /home/ilker/Projects/OpenICEDA/Project/xschem/RingOslHw.sch
**.subckt RingOslHw PD VCTRL VCC VSS VON VOP
*.ipin PD
*.ipin VCTRL
*.iopin VCC
*.iopin VSS
*.opin VON
*.opin VOP
X2 VCC VSS net4 net3 VCTRL PD VOP VON VCC VSS net4 net3 VCTRL PD VOP VON inverterblock
X1 VCC VSS net2 net1 VCTRL PD net3 net4 VCC VSS net2 net1 VCTRL PD net3 net4 inverterblock
X3 VCC VSS VON VOP VCTRL PD net1 net2 VCC VSS VON VOP VCTRL PD net1 net2 inverterblock
**** begin user architecture code

** opencircuitdesign pdks install
.lib /home/ilker/Projects/OpenICEDA/src/open_pdks/sky130/sky130A/libs.tech/ngspice/sky130.lib.spice tt



* this option enables mos model bin
* selection based on W/NF instead of W
.option wnflag=1
*.option savecurrents
.control
tran 0.01n 1us
plot v(VON) vs v(VOP)
plot v(VON) v(VCTRL) (VOP)
op
.endc


**** end user architecture code
**.ends

* expanding   symbol:  inverterblock.sym # of pins=16
** sym_path: /home/ilker/Projects/OpenICEDA/Project/xschem/inverterblock.sym
** sch_path: /home/ilker/Projects/OpenICEDA/Project/xschem/inverterblock.sch
.subckt inverterblock  VCC VSS VON VOP VCTRL PD VIN VIP VCC VSS VON VOP VCTRL PD VIN VIP
*.ipin VIP
*.opin VON
*.opin VOP
*.ipin PD
*.iopin VSS
*.ipin VIN
*.ipin VCTRL
*.iopin VCC
XM9 net1 PD VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM10 VON VCTRL VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 VON VON VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 VON VON VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 VON VCTRL VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 VON VIP net1 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM7 VON VIN net1 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
