** sch_path: /home/ilker/Projects/OpenICEDA/Project/xschem/untitled-1.sch
**.subckt untitled-1 vcc in in vcc vcc out out2
*.opin vcc
*.ipin in
*.ipin in
*.opin vcc
*.opin vcc
*.opin out
*.opin out2
V1 vcc GND 1.8
V2 in GND SIN(0.1 100m 10 0 0)
R1 vcc in 100k m=1
R2 in GND 100k m=1
R4 out2 vcc 1k m=1
XM3 out in out2 out2 sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
R3 out GND 200 m=1
**** begin user architecture code

** opencircuitdesign pdks install
.lib /home/ilker/Projects/OpenICEDA/src/open_pdks/sky130/sky130A/libs.tech/ngspice/sky130.lib.spice tt_mm




.tran 10e-06 100e-03 0e-03
.control
run
plot v(out) v(in) v(out2)
.endc
.end


**** end user architecture code
**.ends
.GLOBAL GND
.end
